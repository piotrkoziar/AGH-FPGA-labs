// Huffman_coder_tb.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module Huffman_coder_tb (
	);

	wire         huffman_coder_inst_clk_bfm_clk_clk;       // Huffman_coder_inst_clk_bfm:clk -> [Huffman_coder_inst:clk_clk, Huffman_coder_inst_exported_out_bfm:clk, Huffman_coder_inst_reset_bfm:clk]
	wire  [31:0] huffman_coder_inst_exported_out_eco;      // Huffman_coder_inst:exported_out_eco -> Huffman_coder_inst_exported_out_bfm:sig_eco
	wire         huffman_coder_inst_exported_out_ebo;      // Huffman_coder_inst:exported_out_ebo -> Huffman_coder_inst_exported_out_bfm:sig_ebo
	wire   [5:0] huffman_coder_inst_exported_out_lno;      // Huffman_coder_inst:exported_out_lno -> Huffman_coder_inst_exported_out_bfm:sig_lno
	wire         huffman_coder_inst_reset_bfm_reset_reset; // Huffman_coder_inst_reset_bfm:reset -> Huffman_coder_inst:reset_reset_n

	Huffman_coder huffman_coder_inst (
		.clk_clk          (huffman_coder_inst_clk_bfm_clk_clk),       //          clk.clk
		.exported_out_ebo (huffman_coder_inst_exported_out_ebo),      // exported_out.ebo
		.exported_out_eco (huffman_coder_inst_exported_out_eco),      //             .eco
		.exported_out_lno (huffman_coder_inst_exported_out_lno),      //             .lno
		.reset_reset_n    (huffman_coder_inst_reset_bfm_reset_reset)  //        reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) huffman_coder_inst_clk_bfm (
		.clk (huffman_coder_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm huffman_coder_inst_exported_out_bfm (
		.clk     (huffman_coder_inst_clk_bfm_clk_clk),  //     clk.clk
		.sig_ebo (huffman_coder_inst_exported_out_ebo), // conduit.ebo
		.sig_eco (huffman_coder_inst_exported_out_eco), //        .eco
		.sig_lno (huffman_coder_inst_exported_out_lno), //        .lno
		.reset   (1'b0)                                 // (terminated)
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) huffman_coder_inst_reset_bfm (
		.reset (huffman_coder_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (huffman_coder_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
